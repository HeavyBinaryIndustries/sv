module RAMSDP
#(bus_width = 8,
	addr_width = 8,
	initfile = "UNUSED",
	device = "Cyclone V")
(input clock,
 input wren,
 input [addr_width-1:0] rdaddress,
 input [addr_width-1:0] wraddress,
 input [bus_width-1:0] data,
 output	logic [bus_width-1:0] q);

	logic [bus_width-1:0] q_ram;
	logic [2:0][bus_width-1:0] data_ff;
        logic [2:0]same_address = 0;

	always_ff @(posedge clock) begin
		data_ff[2] <= data_ff[1];
		data_ff[1] <= data_ff[0];
 		data_ff[0] <= data;
 		same_address <<= 1;
		same_address[0] <= (wraddress == rdaddress) && wren;
 	end

  assign q = same_address[1] ? data_ff[1] : q_ram;

	altsyncram	altsyncram_component (
				.address_a (wraddress),
				.address_b (rdaddress),
				.clock0 (clock),
				.data_a (data),
				.wren_a (wren),
				.q_b (q_ram),
				.aclr0 (1'b0),
				.aclr1 (1'b0),
				.addressstall_a (1'b0),
				.addressstall_b (1'b0),
				.byteena_a (1'b1),
				.byteena_b (1'b1),
				.clock1 (1'b1),
				.clocken0 (1'b1),
				.clocken1 (1'b1),
				.clocken2 (1'b1),
				.clocken3 (1'b1),
				.data_b (0),
				.eccstatus (),
				.q_a (),
				.rden_a (1'b1),
				.rden_b (1'b1),
				.wren_b (1'b0));

	defparam
		altsyncram_component.address_aclr_b = "NONE",
		altsyncram_component.address_reg_b = "CLOCK0",
		altsyncram_component.clock_enable_input_a = "BYPASS",
		altsyncram_component.clock_enable_input_b = "BYPASS",
		altsyncram_component.clock_enable_output_b = "BYPASS",
		altsyncram_component.init_file = initfile,
		altsyncram_component.intended_device_family = device,
		altsyncram_component.lpm_type = "altsyncram",
		altsyncram_component.numwords_a = 2 ** addr_width,
		altsyncram_component.numwords_b = 2 ** addr_width,
		altsyncram_component.operation_mode = "DUAL_PORT",
		altsyncram_component.outdata_aclr_b = "NONE",
		altsyncram_component.outdata_reg_b = "CLOCK0",
		altsyncram_component.power_up_uninitialized = "FALSE",
		altsyncram_component.read_during_write_mode_mixed_ports = "DONT_CARE",
		altsyncram_component.widthad_a = addr_width,
		altsyncram_component.widthad_b = addr_width,
		altsyncram_component.width_a = bus_width,
		altsyncram_component.width_b = bus_width,


altsyncram_component.width_byteena_a = 1;

endmodule
